
//Async 32:5 encoder


module encoder_32(in, out);

	input [31:0] in;
	output reg [4:0] out;
	
	always @(*) begin
	
		     if (in < 32'h00000002) out <= 5'b00000;
		else if (in < 32'h00000004) out <= 5'b00001;
		else if (in < 32'h00000008) out <= 5'b00010;
		else if (in < 32'h00000010) out <= 5'b00011;
		else if (in < 32'h00000020) out <= 5'b00100;
		else if (in < 32'h00000040) out <= 5'b00101;
		else if (in < 32'h00000080) out <= 5'b00110;
		else if (in < 32'h00000100) out <= 5'b00111;
		else if (in < 32'h00000200) out <= 5'b01000;
		else if (in < 32'h00000400) out <= 5'b01001;
		else if (in < 32'h00000800) out <= 5'b01010;
		else if (in < 32'h00001000) out <= 5'b01011;
		else if (in < 32'h00002000) out <= 5'b01100;
		else if (in < 32'h00004000) out <= 5'b01101;
		else if (in < 32'h00008000) out <= 5'b01110;
		else if (in < 32'h00010000) out <= 5'b01111;
		else if (in < 32'h00020000) out <= 5'b10000;
		else if (in < 32'h00040000) out <= 5'b10001;
		else if (in < 32'h00080000) out <= 5'b10010;
		else if (in < 32'h00100000) out <= 5'b10011;
		else if (in < 32'h00200000) out <= 5'b10100;
		else if (in < 32'h00400000) out <= 5'b10101;
		else if (in < 32'h00800000) out <= 5'b10110;
		else if (in < 32'h01000000) out <= 5'b10111;
		else if (in < 32'h02000000) out <= 5'b11000;
		else if (in < 32'h04000000) out <= 5'b11001;
		else if (in < 32'h08000000) out <= 5'b11010;
		else if (in < 32'h10000000) out <= 5'b11011;
		else if (in < 32'h20000000) out <= 5'b11100;
		else if (in < 32'h40000000) out <= 5'b11101;
		else if (in < 32'h80000000) out <= 5'b11110;
		else 								 out <= 5'b11111;
		/*
		case(in)
			32'b00000000000000000000000000000001: out <= 5'b00000;
			32'b00000000000000000000000000000010: out <= 5'b00001;
			32'b00000000000000000000000000000100: out <= 5'b00010;
			32'b00000000000000000000000000001000: out <= 5'b00011;
			32'b00000000000000000000000000010000: out <= 5'b00100;
			32'b00000000000000000000000000100000: out <= 5'b00101;
			32'b00000000000000000000000001000000: out <= 5'b00110;
			32'b00000000000000000000000010000000: out <= 5'b00111;
			32'b00000000000000000000000100000000: out <= 5'b01000;
			32'b00000000000000000000001000000000: out <= 5'b01001;
			32'b00000000000000000000010000000000: out <= 5'b01010;
			32'b00000000000000000000100000000000: out <= 5'b01011;
			32'b00000000000000000001000000000000: out <= 5'b01100;
			32'b00000000000000000010000000000000: out <= 5'b01101;
			32'b00000000000000000100000000000000: out <= 5'b01110;
			32'b00000000000000001000000000000000: out <= 5'b01111;
			32'b00000000000000010000000000000000: out <= 5'b10000;
			32'b00000000000000100000000000000000: out <= 5'b10001;
			32'b00000000000001000000000000000000: out <= 5'b10010;
			32'b00000000000010000000000000000000: out <= 5'b10011;
			32'b00000000000100000000000000000000: out <= 5'b10100;
			32'b00000000001000000000000000000000: out <= 5'b10101;
			32'b00000000010000000000000000000000: out <= 5'b10110;
			32'b00000000100000000000000000000000: out <= 5'b10111;
			32'b00000001000000000000000000000000: out <= 5'b11000;
			32'b00000010000000000000000000000000: out <= 5'b11001;
			32'b00000100000000000000000000000000: out <= 5'b11010;
			32'b00001000000000000000000000000000: out <= 5'b11011;
			32'b00010000000000000000000000000000: out <= 5'b11100;
			32'b00100000000000000000000000000000: out <= 5'b11101;
			32'b01000000000000000000000000000000: out <= 5'b11110;
			32'b10000000000000000000000000000000: out <= 5'b11111;
		endcase
	*/
	end

endmodule